module register_tb;

	/*****************************/
	/* Variables for Input Ports */
	/*****************************/
	reg [31:0] in;
	reg en;
	reg clk;

	/******************************/
	/* Variables for Output Ports */
	/******************************/
	wire [31:0] out;
	
	/*****************/
	/* Instanciation */
	/*****************/
	register r(
		.in(in),
		.out(out),
		.en(en),
		.clk(clk)
	);
	
	/***********/
	/* Initial */
	/***********/
	initial begin
		in = 32'h0000FFFF;
		en = 0;
		clk = 0;
		#1;
		
		in = 32'h0000FFFF;
		en = 0;
		clk = 1;
		#1;
		
		in = 32'h0000FFFF;
		en = 1;
		clk = 0;
		#1;
		
		in = 32'h0000FFFF;
		en = 1;
		clk = 1;
		#1;
	end

endmodule